module slave_top(
    inout SDA,
    input rstn,
    input SCL
);
reg [6:0] slave_addr_reg = 7'b1010101;

acL_TSB tsb0 (.IN               (1'b0),
              .EN               (sda_o),
              .OUT              (SDA)
              );

acH_TSB tsb1 (.IN               (SDA),
              .EN               (sda_in_en),
              .OUT              (sda_i)
              );

tx_fifo fifo (.clk              (SCL),
              .rst              (rstn),
              .wr_en_tx         (wr_en_fifo),
              .rd_en_tx         (rd_en_fifo),
              .data_in          (wr_data),
              .full             (FIFO_FULL),
              .empty            (FIFO_EMPTY),
              .data_out         (rd_data)
              );

clk_div_final div0(.clk_i(clk),
                   .rstn(rstn),
                   .clk_en(clk_en),
                   .clk_s(clk_s),
                   .clk_t(clk_t),
                   .scl(SCL) //assuming the SCL is generated by the clock divider and not an input from the master --> just for debugging
                   );

slave_fsm fsm (.sda_i           (sda_i),
               .clk_t           (clk_t),
               .SCL           (SCL),
               .FIFO_FULL       (FIFO_FULL),
               .FIFO_EMPTY      (FIFO_EMPTY),
               .start_det       (start_det),
               .stop_det        (stop_det),
               .rstn            (rstn),
               .rd_data         (rd_data),
               .slave_addr_reg  (slave_addr_reg),
               .sda_o           (sda_o),
               .sda_in_en       (sda_in_en),
               .wr_en_fifo      (wr_en_fifo),
               .rd_en_fifo      (rd_en_fifo),
               .wr_data         (wr_data)
               );

start_stop_det det (.scl        (clk_s),
                    .sda_i      (SDA),
                    .det_en     (SCL),
                    .rstn       (rstn),
                    .start_det  (start_det),
                    .stop_det   (stop_det)
                    );


endmodule